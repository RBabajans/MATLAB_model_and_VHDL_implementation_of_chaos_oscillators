library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Heaviside_memory is
    Port (
        clk      : in  STD_LOGIC;  -- Clock signal
        we       : in  STD_LOGIC;  -- Write Enable
        addr     : in  STD_LOGIC_VECTOR(11 downto 0); -- 12-bit Address space
        d_in      : in  STD_LOGIC_VECTOR(21 downto 0); -- Data input (22-bit)
        d_out     : out STD_LOGIC_VECTOR(21 downto 0)  -- Data output (22-bit)
    );
end Heaviside_memory;

architecture rtl of Heaviside_memory is

	 signal mem_out_reg, mem_out_next : STD_LOGIC_VECTOR(21 downto 0) := (others => '0');


    type Heaviside_Array is array (0 to 4095) of STD_LOGIC_VECTOR(21 downto 0);  -- Memory array
    signal mem : Heaviside_Array := (
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111111111111111",
"0111111111100000000000",
"0111111110100010000000",
"0111111101100100000000",
"0111111100100110000000",
"0111111011101000000000",
"0111111010101010000000",
"0111111001101100000000",
"0111111000101110000000",
"0111110111110000000000",
"0111110110110010000000",
"0111110101110100000000",
"0111110100110110000000",
"0111110011111000000000",
"0111110010111010000000",
"0111110001111100000000",
"0111110000111110000000",
"0111110000000000000000",
"0111101111000010000000",
"0111101110000100000000",
"0111101101000110000000",
"0111101100001000000000",
"0111101011001010000000",
"0111101010001100000000",
"0111101001001110000000",
"0111101000010000000000",
"0111100111010010000000",
"0111100110010100000000",
"0111100101010110000000",
"0111100100011000000000",
"0111100011011010000000",
"0111100010011100000000",
"0111100001011110000000",
"0111100000100000000000",
"0111011111100010000000",
"0111011110100100000000",
"0111011101100110000000",
"0111011100101000000000",
"0111011011101010000000",
"0111011010101100000000",
"0111011001101110000000",
"0111011000110000000000",
"0111010111110010000000",
"0111010110110100000000",
"0111010101110110000000",
"0111010100111000000000",
"0111010011111010000000",
"0111010010111100000000",
"0111010001111110000000",
"0111010001000000000000",
"0111010000000010000000",
"0111001111000100000000",
"0111001110000110000000",
"0111001101001000000000",
"0111001100001010000000",
"0111001011001100000000",
"0111001010001110000000",
"0111001001010000000000",
"0111001000010010000000",
"0111000111010100000000",
"0111000110010110000000",
"0111000101011000000000",
"0111000100011010000000",
"0111000011011100000000",
"0111000010011110000000",
"0111000001100000000000",
"0111000000100010000000",
"0110111111100100000000",
"0110111110100110000000",
"0110111101101000000000",
"0110111100101010000000",
"0110111011101100000000",
"0110111010101110000000",
"0110111001110000000000",
"0110111000110010000000",
"0110110111110100000000",
"0110110110110110000000",
"0110110101111000000000",
"0110110100111010000000",
"0110110011111100000000",
"0110110010111110000000",
"0110110010000000000000",
"0110110001000010000000",
"0110110000000100000000",
"0110101111000110000000",
"0110101110001000000000",
"0110101101001010000000",
"0110101100001100000000",
"0110101011001110000000",
"0110101010010000000000",
"0110101001010010000000",
"0110101000010100000000",
"0110100111010110000000",
"0110100110011000000000",
"0110100101011010000000",
"0110100100011100000000",
"0110100011011110000000",
"0110100010100000000000",
"0110100001100010000000",
"0110100000100100000000",
"0110011111100110000000",
"0110011110101000000000",
"0110011101101010000000",
"0110011100101100000000",
"0110011011101110000000",
"0110011010110000000000",
"0110011001110010000000",
"0110011000110100000000",
"0110010111110110000000",
"0110010110111000000000",
"0110010101111010000000",
"0110010100111100000000",
"0110010011111110000000",
"0110010011000000000000",
"0110010010000010000000",
"0110010001000100000000",
"0110010000000110000000",
"0110001111001000000000",
"0110001110001010000000",
"0110001101001100000000",
"0110001100001110000000",
"0110001011010000000000",
"0110001010010010000000",
"0110001001010100000000",
"0110001000010110000000",
"0110000111011000000000",
"0110000110011010000000",
"0110000101011100000000",
"0110000100011110000000",
"0110000011100000000000",
"0110000010100010000000",
"0110000001100100000000",
"0110000000100110000000",
"0101111111101000000000",
"0101111110101010000000",
"0101111101101100000000",
"0101111100101110000000",
"0101111011110000000000",
"0101111010110010000000",
"0101111001110100000000",
"0101111000110110000000",
"0101110111111000000000",
"0101110110111010000000",
"0101110101111100000000",
"0101110100111110000000",
"0101110100000000000000",
"0101110011000010000000",
"0101110010000100000000",
"0101110001000110000000",
"0101110000001000000000",
"0101101111001010000000",
"0101101110001100000000",
"0101101101001110000000",
"0101101100010000000000",
"0101101011010010000000",
"0101101010010100000000",
"0101101001010110000000",
"0101101000011000000000",
"0101100111011010000000",
"0101100110011100000000",
"0101100101011110000000",
"0101100100100000000000",
"0101100011100010000000",
"0101100010100100000000",
"0101100001100110000000",
"0101100000101000000000",
"0101011111101010000000",
"0101011110101100000000",
"0101011101101110000000",
"0101011100110000000000",
"0101011011110010000000",
"0101011010110100000000",
"0101011001110110000000",
"0101011000111000000000",
"0101010111111010000000",
"0101010110111100000000",
"0101010101111110000000",
"0101010101000000000000",
"0101010100000010000000",
"0101010011000100000000",
"0101010010000110000000",
"0101010001001000000000",
"0101010000001010000000",
"0101001111001100000000",
"0101001110001110000000",
"0101001101010000000000",
"0101001100010010000000",
"0101001011010100000000",
"0101001010010110000000",
"0101001001011000000000",
"0101001000011010000000",
"0101000111011100000000",
"0101000110011110000000",
"0101000101100000000000",
"0101000100100010000000",
"0101000011100100000000",
"0101000010100110000000",
"0101000001101000000000",
"0101000000101010000000",
"0100111111101100000000",
"0100111110101110000000",
"0100111101110000000000",
"0100111100110010000000",
"0100111011110100000000",
"0100111010110110000000",
"0100111001111000000000",
"0100111000111010000000",
"0100110111111100000000",
"0100110110111110000000",
"0100110110000000000000",
"0100110101000010000000",
"0100110100000100000000",
"0100110011000110000000",
"0100110010001000000000",
"0100110001001010000000",
"0100110000001100000000",
"0100101111001110000000",
"0100101110010000000000",
"0100101101010010000000",
"0100101100010100000000",
"0100101011010110000000",
"0100101010011000000000",
"0100101001011010000000",
"0100101000011100000000",
"0100100111011110000000",
"0100100110100000000000",
"0100100101100010000000",
"0100100100100100000000",
"0100100011100110000000",
"0100100010101000000000",
"0100100001101010000000",
"0100100000101100000000",
"0100011111101110000000",
"0100011110110000000000",
"0100011101110010000000",
"0100011100110100000000",
"0100011011110110000000",
"0100011010111000000000",
"0100011001111010000000",
"0100011000111100000000",
"0100010111111110000000",
"0100010111000000000000",
"0100010110000010000000",
"0100010101000100000000",
"0100010100000110000000",
"0100010011001000000000",
"0100010010001010000000",
"0100010001001100000000",
"0100010000001110000000",
"0100001111010000000000",
"0100001110010010000000",
"0100001101010100000000",
"0100001100010110000000",
"0100001011011000000000",
"0100001010011010000000",
"0100001001011100000000",
"0100001000011110000000",
"0100000111100000000000",
"0100000110100010000000",
"0100000101100100000000",
"0100000100100110000000",
"0100000011101000000000",
"0100000010101010000000",
"0100000001101100000000",
"0100000000101110000000",
"0011111111110000000000",
"0011111110110010000000",
"0011111101110100000000",
"0011111100110110000000",
"0011111011111000000000",
"0011111010111010000000",
"0011111001111100000000",
"0011111000111110000000",
"0011111000000000000000",
"0011110111000010000000",
"0011110110000100000000",
"0011110101000110000000",
"0011110100001000000000",
"0011110011001010000000",
"0011110010001100000000",
"0011110001001110000000",
"0011110000010000000000",
"0011101111010010000000",
"0011101110010100000000",
"0011101101010110000000",
"0011101100011000000000",
"0011101011011010000000",
"0011101010011100000000",
"0011101001011110000000",
"0011101000100000000000",
"0011100111100010000000",
"0011100110100100000000",
"0011100101100110000000",
"0011100100101000000000",
"0011100011101010000000",
"0011100010101100000000",
"0011100001101110000000",
"0011100000110000000000",
"0011011111110010000000",
"0011011110110100000000",
"0011011101110110000000",
"0011011100111000000000",
"0011011011111010000000",
"0011011010111100000000",
"0011011001111110000000",
"0011011001000000000000",
"0011011000000010000000",
"0011010111000100000000",
"0011010110000110000000",
"0011010101001000000000",
"0011010100001010000000",
"0011010011001100000000",
"0011010010001110000000",
"0011010001010000000000",
"0011010000010010000000",
"0011001111010100000000",
"0011001110010110000000",
"0011001101011000000000",
"0011001100011010000000",
"0011001011011100000000",
"0011001010011110000000",
"0011001001100000000000",
"0011001000100010000000",
"0011000111100100000000",
"0011000110100110000000",
"0011000101101000000000",
"0011000100101010000000",
"0011000011101100000000",
"0011000010101110000000",
"0011000001110000000000",
"0011000000110010000000",
"0010111111110100000000",
"0010111110110110000000",
"0010111101111000000000",
"0010111100111010000000",
"0010111011111100000000",
"0010111010111110000000",
"0010111010000000000000",
"0010111001000010000000",
"0010111000000100000000",
"0010110111000110000000",
"0010110110001000000000",
"0010110101001010000000",
"0010110100001100000000",
"0010110011001110000000",
"0010110010010000000000",
"0010110001010010000000",
"0010110000010100000000",
"0010101111010110000000",
"0010101110011000000000",
"0010101101011010000000",
"0010101100011100000000",
"0010101011011110000000",
"0010101010100000000000",
"0010101001100010000000",
"0010101000100100000000",
"0010100111100110000000",
"0010100110101000000000",
"0010100101101010000000",
"0010100100101100000000",
"0010100011101110000000",
"0010100010110000000000",
"0010100001110010000000",
"0010100000110100000000",
"0010011111110110000000",
"0010011110111000000000",
"0010011101111010000000",
"0010011100111100000000",
"0010011011111110000000",
"0010011011000000000000",
"0010011010000010000000",
"0010011001000100000000",
"0010011000000110000000",
"0010010111001000000000",
"0010010110001010000000",
"0010010101001100000000",
"0010010100001110000000",
"0010010011010000000000",
"0010010010010010000000",
"0010010001010100000000",
"0010010000010110000000",
"0010001111011000000000",
"0010001110011010000000",
"0010001101011100000000",
"0010001100011110000000",
"0010001011100000000000",
"0010001010100010000000",
"0010001001100100000000",
"0010001000100110000000",
"0010000111101000000000",
"0010000110101010000000",
"0010000101101100000000",
"0010000100101110000000",
"0010000011110000000000",
"0010000010110010000000",
"0010000001110100000000",
"0010000000110110000000",
"0001111111111000000000",
"0001111110111010000000",
"0001111101111100000000",
"0001111100111110000000",
"0001111100000000000000",
"0001111011000010000000",
"0001111010000100000000",
"0001111001000110000000",
"0001111000001000000000",
"0001110111001010000000",
"0001110110001100000000",
"0001110101001110000000",
"0001110100010000000000",
"0001110011010010000000",
"0001110010010100000000",
"0001110001010110000000",
"0001110000011000000000",
"0001101111011010000000",
"0001101110011100000000",
"0001101101011110000000",
"0001101100100000000000",
"0001101011100010000000",
"0001101010100100000000",
"0001101001100110000000",
"0001101000101000000000",
"0001100111101010000000",
"0001100110101100000000",
"0001100101101110000000",
"0001100100110000000000",
"0001100011110010000000",
"0001100010110100000000",
"0001100001110110000000",
"0001100000111000000000",
"0001011111111010000000",
"0001011110111100000000",
"0001011101111110000000",
"0001011101000000000000",
"0001011100000010000000",
"0001011011000100000000",
"0001011010000110000000",
"0001011001001000000000",
"0001011000001010000000",
"0001010111001100000000",
"0001010110001110000000",
"0001010101010000000000",
"0001010100010010000000",
"0001010011010100000000",
"0001010010010110000000",
"0001010001011000000000",
"0001010000011010000000",
"0001001111011100000000",
"0001001110011110000000",
"0001001101100000000000",
"0001001100100010000000",
"0001001011100100000000",
"0001001010100110000000",
"0001001001101000000000",
"0001001000101010000000",
"0001000111101100000000",
"0001000110101110000000",
"0001000101110000000000",
"0001000100110010000000",
"0001000011110100000000",
"0001000010110110000000",
"0001000001111000000000",
"0001000000111010000000",
"0000111111111100000000",
"0000111110111110000000",
"0000111110000000000000",
"0000111101000010000000",
"0000111100000100000000",
"0000111011000110000000",
"0000111010001000000000",
"0000111001001010000000",
"0000111000001100000000",
"0000110111001110000000",
"0000110110010000000000",
"0000110101010010000000",
"0000110100010100000000",
"0000110011010110000000",
"0000110010011000000000",
"0000110001011010000000",
"0000110000011100000000",
"0000101111011110000000",
"0000101110100000000000",
"0000101101100010000000",
"0000101100100100000000",
"0000101011100110000000",
"0000101010101000000000",
"0000101001101010000000",
"0000101000101100000000",
"0000100111101110000000",
"0000100110110000000000",
"0000100101110010000000",
"0000100100110100000000",
"0000100011110110000000",
"0000100010111000000000",
"0000100001111010000000",
"0000100000111100000000",
"0000011111111110000000",
"0000011111000000000000",
"0000011110000010000000",
"0000011101000100000000",
"0000011100000110000000",
"0000011011001000000000",
"0000011010001010000000",
"0000011001001100000000",
"0000011000001110000000",
"0000010111010000000000",
"0000010110010010000000",
"0000010101010100000000",
"0000010100010110000000",
"0000010011011000000000",
"0000010010011010000000",
"0000010001011100000000",
"0000010000011110000000",
"0000001111100000000000",
"0000001110100010000000",
"0000001101100100000000",
"0000001100100110000000",
"0000001011101000000000",
"0000001010101010000000",
"0000001001101100000000",
"0000001000101110000000",
"0000000111110000000000",
"0000000110110010000000",
"0000000101110100000000",
"0000000100110110000000",
"0000000011111000000000",
"0000000010111010000000",
"0000000001111100000000",
"0000000000111110000000",
"0000000000000000000000",
"1111111111000010000000",
"1111111110000100000000",
"1111111101000110000000",
"1111111100001000000000",
"1111111011001010000000",
"1111111010001100000000",
"1111111001001110000000",
"1111111000010000000000",
"1111110111010010000000",
"1111110110010100000000",
"1111110101010110000000",
"1111110100011000000000",
"1111110011011010000000",
"1111110010011100000000",
"1111110001011110000000",
"1111110000100000000000",
"1111101111100010000000",
"1111101110100100000000",
"1111101101100110000000",
"1111101100101000000000",
"1111101011101010000000",
"1111101010101100000000",
"1111101001101110000000",
"1111101000110000000000",
"1111100111110010000000",
"1111100110110100000000",
"1111100101110110000000",
"1111100100111000000000",
"1111100011111010000000",
"1111100010111100000000",
"1111100001111110000000",
"1111100001000000000000",
"1111100000000010000000",
"1111011111000100000000",
"1111011110000110000000",
"1111011101001000000000",
"1111011100001010000000",
"1111011011001100000000",
"1111011010001110000000",
"1111011001010000000000",
"1111011000010010000000",
"1111010111010100000000",
"1111010110010110000000",
"1111010101011000000000",
"1111010100011010000000",
"1111010011011100000000",
"1111010010011110000000",
"1111010001100000000000",
"1111010000100010000000",
"1111001111100100000000",
"1111001110100110000000",
"1111001101101000000000",
"1111001100101010000000",
"1111001011101100000000",
"1111001010101110000000",
"1111001001110000000000",
"1111001000110010000000",
"1111000111110100000000",
"1111000110110110000000",
"1111000101111000000000",
"1111000100111010000000",
"1111000011111100000000",
"1111000010111110000000",
"1111000010000000000000",
"1111000001111010011010",
"1111000001110100110101",
"1111000001101111001111",
"1111000001101001101001",
"1111000001100100000011",
"1111000001011110011110",
"1111000001011000111000",
"1111000001010011010010",
"1111000001001101101100",
"1111000001001000000111",
"1111000001000010100001",
"1111000000111100111011",
"1111000000110111010101",
"1111000000110001110000",
"1111000000101100001010",
"1111000000100110100100",
"1111000000100000111110",
"1111000000011011011001",
"1111000000010101110011",
"1111000000010000001101",
"1111000000001010100111",
"1111000000000101000010",
"1110111111111111011100",
"1110111111111001110110",
"1110111111110100010000",
"1110111111101110101011",
"1110111111101001000101",
"1110111111100011011111",
"1110111111011101111001",
"1110111111011000010100",
"1110111111010010101110",
"1110111111001101001000",
"1110111111000111100010",
"1110111111000001111101",
"1110111110111100010111",
"1110111110110110110001",
"1110111110110001001011",
"1110111110101011100110",
"1110111110100110000000",
"1110111110100000011010",
"1110111110011010110101",
"1110111110010101001111",
"1110111110001111101001",
"1110111110001010000011",
"1110111110000100011110",
"1110111101111110111000",
"1110111101111001010010",
"1110111101110011101100",
"1110111101101110000111",
"1110111101101000100001",
"1110111101100010111011",
"1110111101011101010101",
"1110111101010111110000",
"1110111101010010001010",
"1110111101001100100100",
"1110111101000110111110",
"1110111101000001011001",
"1110111100111011110011",
"1110111100110110001101",
"1110111100110000100111",
"1110111100101011000010",
"1110111100100101011100",
"1110111100011111110110",
"1110111100011010010000",
"1110111100010100101011",
"1110111100001111000101",
"1110111100001001011111",
"1110111100000011111001",
"1110111011111110010100",
"1110111011111000101110",
"1110111011110011001000",
"1110111011101101100010",
"1110111011100111111101",
"1110111011100010010111",
"1110111011011100110001",
"1110111011010111001011",
"1110111011010001100110",
"1110111011001100000000",
"1110111011000110011010",
"1110111011000000110101",
"1110111010111011001111",
"1110111010110101101001",
"1110111010110000000011",
"1110111010101010011110",
"1110111010100100111000",
"1110111010011111010010",
"1110111010011001101100",
"1110111010010100000111",
"1110111010001110100001",
"1110111010001000111011",
"1110111010000011010101",
"1110111001111101110000",
"1110111001111000001010",
"1110111001110010100100",
"1110111001101100111110",
"1110111001100111011001",
"1110111001100001110011",
"1110111001011100001101",
"1110111001010110100111",
"1110111001010001000010",
"1110111001001011011100",
"1110111001000101110110",
"1110111001000000010000",
"1110111000111010101011",
"1110111000110101000101",
"1110111000101111011111",
"1110111000101001111001",
"1110111000100100010100",
"1110111000011110101110",
"1110111000011001001000",
"1110111000010011100010",
"1110111000001101111101",
"1110111000001000010111",
"1110111000000010110001",
"1110110111111101001011",
"1110110111110111100110",
"1110110111110010000000",
"1110110111101100011010",
"1110110111100110110101",
"1110110111100001001111",
"1110110111011011101001",
"1110110111010110000011",
"1110110111010000011110",
"1110110111001010111000",
"1110110111000101010010",
"1110110110111111101100",
"1110110110111010000111",
"1110110110110100100001",
"1110110110101110111011",
"1110110110101001010101",
"1110110110100011110000",
"1110110110011110001010",
"1110110110011000100100",
"1110110110010010111110",
"1110110110001101011001",
"1110110110000111110011",
"1110110110000010001101",
"1110110101111100100111",
"1110110101110111000010",
"1110110101110001011100",
"1110110101101011110110",
"1110110101100110010000",
"1110110101100000101011",
"1110110101011011000101",
"1110110101010101011111",
"1110110101001111111001",
"1110110101001010010100",
"1110110101000100101110",
"1110110100111111001000",
"1110110100111001100010",
"1110110100110011111101",
"1110110100101110010111",
"1110110100101000110001",
"1110110100100011001011",
"1110110100011101100110",
"1110110100011000000000",
"1110110100010010011010",
"1110110100001100110101",
"1110110100000111001111",
"1110110100000001101001",
"1110110011111100000011",
"1110110011110110011110",
"1110110011110000111000",
"1110110011101011010010",
"1110110011100101101100",
"1110110011100000000111",
"1110110011011010100001",
"1110110011010100111011",
"1110110011001111010101",
"1110110011001001110000",
"1110110011000100001010",
"1110110010111110100100",
"1110110010111000111110",
"1110110010110011011001",
"1110110010101101110011",
"1110110010101000001101",
"1110110010100010100111",
"1110110010011101000010",
"1110110010010111011100",
"1110110010010001110110",
"1110110010001100010000",
"1110110010000110101011",
"1110110010000001000101",
"1110110001111011011111",
"1110110001110101111001",
"1110110001110000010100",
"1110110001101010101110",
"1110110001100101001000",
"1110110001011111100010",
"1110110001011001111101",
"1110110001010100010111",
"1110110001001110110001",
"1110110001001001001011",
"1110110001000011100110",
"1110110000111110000000",
"1110110000111000011010",
"1110110000110010110101",
"1110110000101101001111",
"1110110000100111101001",
"1110110000100010000011",
"1110110000011100011110",
"1110110000010110111000",
"1110110000010001010010",
"1110110000001011101100",
"1110110000000110000111",
"1110110000000000100001",
"1110101111111010111011",
"1110101111110101010101",
"1110101111101111110000",
"1110101111101010001010",
"1110101111100100100100",
"1110101111011110111110",
"1110101111011001011001",
"1110101111010011110011",
"1110101111001110001101",
"1110101111001000100111",
"1110101111000011000010",
"1110101110111101011100",
"1110101110110111110110",
"1110101110110010010000",
"1110101110101100101011",
"1110101110100111000101",
"1110101110100001011111",
"1110101110011011111001",
"1110101110010110010100",
"1110101110010000101110",
"1110101110001011001000",
"1110101110000101100010",
"1110101101111111111101",
"1110101101111010010111",
"1110101101110100110001",
"1110101101101111001011",
"1110101101101001100110",
"1110101101100100000000",
"1110101101011110011010",
"1110101101011000110101",
"1110101101010011001111",
"1110101101001101101001",
"1110101101001000000011",
"1110101101000010011110",
"1110101100111100111000",
"1110101100110111010010",
"1110101100110001101100",
"1110101100101100000111",
"1110101100100110100001",
"1110101100100000111011",
"1110101100011011010101",
"1110101100010101110000",
"1110101100010000001010",
"1110101100001010100100",
"1110101100000100111110",
"1110101011111111011001",
"1110101011111001110011",
"1110101011110100001101",
"1110101011101110100111",
"1110101011101001000010",
"1110101011100011011100",
"1110101011011101110110",
"1110101011011000010000",
"1110101011010010101011",
"1110101011001101000101",
"1110101011000111011111",
"1110101011000001111001",
"1110101010111100010100",
"1110101010110110101110",
"1110101010110001001000",
"1110101010101011100010",
"1110101010100101111101",
"1110101010100000010111",
"1110101010011010110001",
"1110101010010101001011",
"1110101010001111100110",
"1110101010001010000000",
"1110101010000100011010",
"1110101001111110110101",
"1110101001111001001111",
"1110101001110011101001",
"1110101001101110000011",
"1110101001101000011110",
"1110101001100010111000",
"1110101001011101010010",
"1110101001010111101100",
"1110101001010010000111",
"1110101001001100100001",
"1110101001000110111011",
"1110101001000001010101",
"1110101000111011110000",
"1110101000110110001010",
"1110101000110000100100",
"1110101000101010111110",
"1110101000100101011001",
"1110101000011111110011",
"1110101000011010001101",
"1110101000010100100111",
"1110101000001111000010",
"1110101000001001011100",
"1110101000000011110110",
"1110100111111110010000",
"1110100111111000101011",
"1110100111110011000101",
"1110100111101101011111",
"1110100111100111111001",
"1110100111100010010100",
"1110100111011100101110",
"1110100111010111001000",
"1110100111010001100010",
"1110100111001011111101",
"1110100111000110010111",
"1110100111000000110001",
"1110100110111011001011",
"1110100110110101100110",
"1110100110110000000000",
"1110100110101010011010",
"1110100110100100110101",
"1110100110011111001111",
"1110100110011001101001",
"1110100110010100000011",
"1110100110001110011110",
"1110100110001000111000",
"1110100110000011010010",
"1110100101111101101100",
"1110100101111000000111",
"1110100101110010100001",
"1110100101101100111011",
"1110100101100111010101",
"1110100101100001110000",
"1110100101011100001010",
"1110100101010110100100",
"1110100101010000111110",
"1110100101001011011001",
"1110100101000101110011",
"1110100101000000001101",
"1110100100111010100111",
"1110100100110101000010",
"1110100100101111011100",
"1110100100101001110110",
"1110100100100100010000",
"1110100100011110101011",
"1110100100011001000101",
"1110100100010011011111",
"1110100100001101111001",
"1110100100001000010100",
"1110100100000010101110",
"1110100011111101001000",
"1110100011110111100010",
"1110100011110001111101",
"1110100011101100010111",
"1110100011100110110001",
"1110100011100001001011",
"1110100011011011100110",
"1110100011010110000000",
"1110100011010000011010",
"1110100011001010110101",
"1110100011000101001111",
"1110100010111111101001",
"1110100010111010000011",
"1110100010110100011110",
"1110100010101110111000",
"1110100010101001010010",
"1110100010100011101100",
"1110100010011110000111",
"1110100010011000100001",
"1110100010010010111011",
"1110100010001101010101",
"1110100010000111110000",
"1110100010000010001010",
"1110100001111100100100",
"1110100001110110111110",
"1110100001110001011001",
"1110100001101011110011",
"1110100001100110001101",
"1110100001100000100111",
"1110100001011011000010",
"1110100001010101011100",
"1110100001001111110110",
"1110100001001010010000",
"1110100001000100101011",
"1110100000111111000101",
"1110100000111001011111",
"1110100000110011111001",
"1110100000101110010100",
"1110100000101000101110",
"1110100000100011001000",
"1110100000011101100010",
"1110100000010111111101",
"1110100000010010010111",
"1110100000001100110001",
"1110100000000111001011",
"1110100000000001100110",
"1110011111111100000000",
"1110011111110110011010",
"1110011111110000110101",
"1110011111101011001111",
"1110011111100101101001",
"1110011111100000000011",
"1110011111011010011110",
"1110011111010100111000",
"1110011111001111010010",
"1110011111001001101100",
"1110011111000100000111",
"1110011110111110100001",
"1110011110111000111011",
"1110011110110011010101",
"1110011110101101110000",
"1110011110101000001010",
"1110011110100010100100",
"1110011110011100111110",
"1110011110010111011001",
"1110011110010001110011",
"1110011110001100001101",
"1110011110000110100111",
"1110011110000001000010",
"1110011101111011011100",
"1110011101110101110110",
"1110011101110000010000",
"1110011101101010101011",
"1110011101100101000101",
"1110011101011111011111",
"1110011101011001111001",
"1110011101010100010100",
"1110011101001110101110",
"1110011101001001001000",
"1110011101000011100010",
"1110011100111101111101",
"1110011100111000010111",
"1110011100110010110001",
"1110011100101101001011",
"1110011100100111100110",
"1110011100100010000000",
"1110011100011100011010",
"1110011100010110110101",
"1110011100010001001111",
"1110011100001011101001",
"1110011100000110000011",
"1110011100000000011110",
"1110011011111010111000",
"1110011011110101010010",
"1110011011101111101100",
"1110011011101010000111",
"1110011011100100100001",
"1110011011011110111011",
"1110011011011001010101",
"1110011011010011110000",
"1110011011001110001010",
"1110011011001000100100",
"1110011011000010111110",
"1110011010111101011001",
"1110011010110111110011",
"1110011010110010001101",
"1110011010101100100111",
"1110011010100111000010",
"1110011010100001011100",
"1110011010011011110110",
"1110011010010110010000",
"1110011010010000101011",
"1110011010001011000101",
"1110011010000101011111",
"1110011001111111111001",
"1110011001111010010100",
"1110011001110100101110",
"1110011001101111001000",
"1110011001101001100010",
"1110011001100011111101",
"1110011001011110010111",
"1110011001011000110001",
"1110011001010011001011",
"1110011001001101100110",
"1110011001001000000000",
"1110011001000010011010",
"1110011000111100110101",
"1110011000110111001111",
"1110011000110001101001",
"1110011000101100000011",
"1110011000100110011110",
"1110011000100000111000",
"1110011000011011010010",
"1110011000010101101100",
"1110011000010000000111",
"1110011000001010100001",
"1110011000000100111011",
"1110010111111111010101",
"1110010111111001110000",
"1110010111110100001010",
"1110010111101110100100",
"1110010111101000111110",
"1110010111100011011001",
"1110010111011101110011",
"1110010111011000001101",
"1110010111010010100111",
"1110010111001101000010",
"1110010111000111011100",
"1110010111000001110110",
"1110010110111100010000",
"1110010110110110101011",
"1110010110110001000101",
"1110010110101011011111",
"1110010110100101111001",
"1110010110100000010100",
"1110010110011010101110",
"1110010110010101001000",
"1110010110001111100010",
"1110010110001001111101",
"1110010110000100010111",
"1110010101111110110001",
"1110010101111001001011",
"1110010101110011100110",
"1110010101101110000000",
"1110010101101000011010",
"1110010101100010110101",
"1110010101011101001111",
"1110010101010111101001",
"1110010101010010000011",
"1110010101001100011110",
"1110010101000110111000",
"1110010101000001010010",
"1110010100111011101100",
"1110010100110110000111",
"1110010100110000100001",
"1110010100101010111011",
"1110010100100101010101",
"1110010100011111110000",
"1110010100011010001010",
"1110010100010100100100",
"1110010100001110111110",
"1110010100001001011001",
"1110010100000011110011",
"1110010011111110001101",
"1110010011111000100111",
"1110010011110011000010",
"1110010011101101011100",
"1110010011100111110110",
"1110010011100010010000",
"1110010011011100101011",
"1110010011010111000101",
"1110010011010001011111",
"1110010011001011111001",
"1110010011000110010100",
"1110010011000000101110",
"1110010010111011001000",
"1110010010110101100010",
"1110010010101111111101",
"1110010010101010010111",
"1110010010100100110001",
"1110010010011111001011",
"1110010010011001100110",
"1110010010010100000000",
"1110010010001110011010",
"1110010010001000110101",
"1110010010000011001111",
"1110010001111101101001",
"1110010001111000000011",
"1110010001110010011110",
"1110010001101100111000",
"1110010001100111010010",
"1110010001100001101100",
"1110010001011100000111",
"1110010001010110100001",
"1110010001010000111011",
"1110010001001011010101",
"1110010001000101110000",
"1110010001000000001010",
"1110010000111010100100",
"1110010000110100111110",
"1110010000101111011001",
"1110010000101001110011",
"1110010000100100001101",
"1110010000011110100111",
"1110010000011001000010",
"1110010000010011011100",
"1110010000001101110110",
"1110010000001000010000",
"1110010000000010101011",
"1110001111111101000101",
"1110001111110111011111",
"1110001111110001111001",
"1110001111101100010100",
"1110001111100110101110",
"1110001111100001001000",
"1110001111011011100010",
"1110001111010101111101",
"1110001111010000010111",
"1110001111001010110001",
"1110001111000101001011",
"1110001110111111100110",
"1110001110111010000000",
"1110001110110100011010",
"1110001110101110110101",
"1110001110101001001111",
"1110001110100011101001",
"1110001110011110000011",
"1110001110011000011110",
"1110001110010010111000",
"1110001110001101010010",
"1110001110000111101100",
"1110001110000010000111",
"1110001101111100100001",
"1110001101110110111011",
"1110001101110001010101",
"1110001101101011110000",
"1110001101100110001010",
"1110001101100000100100",
"1110001101011010111110",
"1110001101010101011001",
"1110001101001111110011",
"1110001101001010001101",
"1110001101000100100111",
"1110001100111111000010",
"1110001100111001011100",
"1110001100110011110110",
"1110001100101110010000",
"1110001100101000101011",
"1110001100100011000101",
"1110001100011101011111",
"1110001100010111111001",
"1110001100010010010100",
"1110001100001100101110",
"1110001100000111001000",
"1110001100000001100010",
"1110001011111011111101",
"1110001011110110010111",
"1110001011110000110001",
"1110001011101011001011",
"1110001011100101100110",
"1110001011100000000000",
"1110001011011010011010",
"1110001011010100110101",
"1110001011001111001111",
"1110001011001001101001",
"1110001011000100000011",
"1110001010111110011110",
"1110001010111000111000",
"1110001010110011010010",
"1110001010101101101100",
"1110001010101000000111",
"1110001010100010100001",
"1110001010011100111011",
"1110001010010111010101",
"1110001010010001110000",
"1110001010001100001010",
"1110001010000110100100",
"1110001010000000111110",
"1110001001111011011001",
"1110001001110101110011",
"1110001001110000001101",
"1110001001101010100111",
"1110001001100101000010",
"1110001001011111011100",
"1110001001011001110110",
"1110001001010100010000",
"1110001001001110101011",
"1110001001001001000101",
"1110001001000011011111",
"1110001000111101111001",
"1110001000111000010100",
"1110001000110010101110",
"1110001000101101001000",
"1110001000100111100010",
"1110001000100001111101",
"1110001000011100010111",
"1110001000010110110001",
"1110001000010001001011",
"1110001000001011100110",
"1110001000000110000000",
"1110001000000000011010",
"1110000111111010110101",
"1110000111110101001111",
"1110000111101111101001",
"1110000111101010000011",
"1110000111100100011110",
"1110000111011110111000",
"1110000111011001010010",
"1110000111010011101100",
"1110000111001110000111",
"1110000111001000100001",
"1110000111000010111011",
"1110000110111101010101",
"1110000110110111110000",
"1110000110110010001010",
"1110000110101100100100",
"1110000110100110111110",
"1110000110100001011001",
"1110000110011011110011",
"1110000110010110001101",
"1110000110010000100111",
"1110000110001011000010",
"1110000110000101011100",
"1110000101111111110110",
"1110000101111010010000",
"1110000101110100101011",
"1110000101101111000101",
"1110000101101001011111",
"1110000101100011111001",
"1110000101011110010100",
"1110000101011000101110",
"1110000101010011001000",
"1110000101001101100010",
"1110000101000111111101",
"1110000101000010010111",
"1110000100111100110001",
"1110000100110111001011",
"1110000100110001100110",
"1110000100101100000000",
"1110000100100110011010",
"1110000100100000110101",
"1110000100011011001111",
"1110000100010101101001",
"1110000100010000000011",
"1110000100001010011110",
"1110000100000100111000",
"1110000011111111010010",
"1110000011111001101100",
"1110000011110100000111",
"1110000011101110100001",
"1110000011101000111011",
"1110000011100011010101",
"1110000011011101110000",
"1110000011011000001010",
"1110000011010010100100",
"1110000011001100111110",
"1110000011000111011001",
"1110000011000001110011",
"1110000010111100001101",
"1110000010110110100111",
"1110000010110001000010",
"1110000010101011011100",
"1110000010100101110110",
"1110000010100000010000",
"1110000010011010101011",
"1110000010010101000101",
"1110000010001111011111",
"1110000010001001111001",
"1110000010000100010100",
"1110000001111110101110",
"1110000001111001001000",
"1110000001110011100010",
"1110000001101101111101",
"1110000001101000010111",
"1110000001100010110001",
"1110000001011101001011",
"1110000001010111100110",
"1110000001010010000000",
"1110000001001100011010",
"1110000001000110110101",
"1110000001000001001111",
"1110000000111011101001",
"1110000000110110000011",
"1110000000110000011110",
"1110000000101010111000",
"1110000000100101010010",
"1110000000011111101100",
"1110000000011010000111",
"1110000000010100100001",
"1110000000001110111011",
"1110000000001001010101",
"1110000000000011110000",
"1101111111111110001010",
"1101111111111000100100",
"1101111111110010111110",
"1101111111101101011001",
"1101111111100111110011",
"1101111111100010001101",
"1101111111011100100111",
"1101111111010111000010",
"1101111111010001011100",
"1101111111001011110110",
"1101111111000110010000",
"1101111111000000101011",
"1101111110111011000101",
"1101111110110101011111",
"1101111110101111111001",
"1101111110101010010100",
"1101111110100100101110",
"1101111110011111001000",
"1101111110011001100010",
"1101111110010011111101",
"1101111110001110010111",
"1101111110001000110001",
"1101111110000011001011",
"1101111101111101100110",
"1101111101111000000000",
"1101111101110010011010",
"1101111101101100110101",
"1101111101100111001111",
"1101111101100001101001",
"1101111101011100000011",
"1101111101010110011110",
"1101111101010000111000",
"1101111101001011010010",
"1101111101000101101100",
"1101111101000000000111",
"1101111100111010100001",
"1101111100110100111011",
"1101111100101111010101",
"1101111100101001110000",
"1101111100100100001010",
"1101111100011110100100",
"1101111100011000111110",
"1101111100010011011001",
"1101111100001101110011",
"1101111100001000001101",
"1101111100000010100111",
"1101111011111101000010",
"1101111011110111011100",
"1101111011110001110110",
"1101111011101100010000",
"1101111011100110101011",
"1101111011100001000101",
"1101111011011011011111",
"1101111011010101111001",
"1101111011010000010100",
"1101111011001010101110",
"1101111011000101001000",
"1101111010111111100010",
"1101111010111001111101",
"1101111010110100010111",
"1101111010101110110001",
"1101111010101001001011",
"1101111010100011100110",
"1101111010011110000000",
"1101111010011000011010",
"1101111010010010110101",
"1101111010001101001111",
"1101111010000111101001",
"1101111010000010000011",
"1101111001111100011110",
"1101111001110110111000",
"1101111001110001010010",
"1101111001101011101100",
"1101111001100110000111",
"1101111001100000100001",
"1101111001011010111011",
"1101111001010101010101",
"1101111001001111110000",
"1101111001001010001010",
"1101111001000100100100",
"1101111000111110111110",
"1101111000111001011001",
"1101111000110011110011",
"1101111000101110001101",
"1101111000101000100111",
"1101111000100011000010",
"1101111000011101011100",
"1101111000010111110110",
"1101111000010010010000",
"1101111000001100101011",
"1101111000000111000101",
"1101111000000001011111",
"1101110111111011111001",
"1101110111110110010100",
"1101110111110000101110",
"1101110111101011001000",
"1101110111100101100010",
"1101110111011111111101",
"1101110111011010010111",
"1101110111010100110001",
"1101110111001111001011",
"1101110111001001100110",
"1101110111000100000000",
"1101110110111110011010",
"1101110110111000110101",
"1101110110110011001111",
"1101110110101101101001",
"1101110110101000000011",
"1101110110100010011110",
"1101110110011100111000",
"1101110110010111010010",
"1101110110010001101100",
"1101110110001100000111",
"1101110110000110100001",
"1101110110000000111011",
"1101110101111011010101",
"1101110101110101110000",
"1101110101110000001010",
"1101110101101010100100",
"1101110101100100111110",
"1101110101011111011001",
"1101110101011001110011",
"1101110101010100001101",
"1101110101001110100111",
"1101110101001001000010",
"1101110101000011011100",
"1101110100111101110110",
"1101110100111000010000",
"1101110100110010101011",
"1101110100101101000101",
"1101110100100111011111",
"1101110100100001111001",
"1101110100011100010100",
"1101110100010110101110",
"1101110100010001001000",
"1101110100001011100010",
"1101110100000101111101",
"1101110100000000010111",
"1101110011111010110001",
"1101110011110101001011",
"1101110011101111100110",
"1101110011101010000000",
"1101110011100100011010",
"1101110011011110110101",
"1101110011011001001111",
"1101110011010011101001",
"1101110011001110000011",
"1101110011001000011110",
"1101110011000010111000",
"1101110010111101010010",
"1101110010110111101100",
"1101110010110010000111",
"1101110010101100100001",
"1101110010100110111011",
"1101110010100001010101",
"1101110010011011110000",
"1101110010010110001010",
"1101110010010000100100",
"1101110010001010111110",
"1101110010000101011001",
"1101110001111111110011",
"1101110001111010001101",
"1101110001110100100111",
"1101110001101111000010",
"1101110001101001011100",
"1101110001100011110110",
"1101110001011110010000",
"1101110001011000101011",
"1101110001010011000101",
"1101110001001101011111",
"1101110001000111111001",
"1101110001000010010100",
"1101110000111100101110",
"1101110000110111001000",
"1101110000110001100010",
"1101110000101011111101",
"1101110000100110010111",
"1101110000100000110001",
"1101110000011011001011",
"1101110000010101100110",
"1101110000010000000000",
"1101110000001010011010",
"1101110000000100110101",
"1101101111111111001111",
"1101101111111001101001",
"1101101111110100000011",
"1101101111101110011110",
"1101101111101000111000",
"1101101111100011010010",
"1101101111011101101100",
"1101101111011000000111",
"1101101111010010100001",
"1101101111001100111011",
"1101101111000111010101",
"1101101111000001110000",
"1101101110111100001010",
"1101101110110110100100",
"1101101110110000111110",
"1101101110101011011001",
"1101101110100101110011",
"1101101110100000001101",
"1101101110011010100111",
"1101101110010101000010",
"1101101110001111011100",
"1101101110001001110110",
"1101101110000100010000",
"1101101101111110101011",
"1101101101111001000101",
"1101101101110011011111",
"1101101101101101111001",
"1101101101101000010100",
"1101101101100010101110",
"1101101101011101001000",
"1101101101010111100010",
"1101101101010001111101",
"1101101101001100010111",
"1101101101000110110001",
"1101101101000001001011",
"1101101100111011100110",
"1101101100110110000000",
"1101101100110000011010",
"1101101100101010110101",
"1101101100100101001111",
"1101101100011111101001",
"1101101100011010000011",
"1101101100010100011110",
"1101101100001110111000",
"1101101100001001010010",
"1101101100000011101100",
"1101101011111110000111",
"1101101011111000100001",
"1101101011110010111011",
"1101101011101101010101",
"1101101011100111110000",
"1101101011100010001010",
"1101101011011100100100",
"1101101011010110111110",
"1101101011010001011001",
"1101101011001011110011",
"1101101011000110001101",
"1101101011000000100111",
"1101101010111011000010",
"1101101010110101011100",
"1101101010101111110110",
"1101101010101010010000",
"1101101010100100101011",
"1101101010011111000101",
"1101101010011001011111",
"1101101010010011111001",
"1101101010001110010100",
"1101101010001000101110",
"1101101010000011001000",
"1101101001111101100010",
"1101101001110111111101",
"1101101001110010010111",
"1101101001101100110001",
"1101101001100111001011",
"1101101001100001100110",
"1101101001011100000000",
"1101101001010110011010",
"1101101001010000110101",
"1101101001001011001111",
"1101101001000101101001",
"1101101001000000000011",
"1101101000111010011110",
"1101101000110100111000",
"1101101000101111010010",
"1101101000101001101100",
"1101101000100100000111",
"1101101000011110100001",
"1101101000011000111011",
"1101101000010011010101",
"1101101000001101110000",
"1101101000001000001010",
"1101101000000010100100",
"1101100111111100111110",
"1101100111110111011001",
"1101100111110001110011",
"1101100111101100001101",
"1101100111100110100111",
"1101100111100001000010",
"1101100111011011011100",
"1101100111010101110110",
"1101100111010000010000",
"1101100111001010101011",
"1101100111000101000101",
"1101100110111111011111",
"1101100110111001111001",
"1101100110110100010100",
"1101100110101110101110",
"1101100110101001001000",
"1101100110100011100010",
"1101100110011101111101",
"1101100110011000010111",
"1101100110010010110001",
"1101100110001101001011",
"1101100110000111100110",
"1101100110000010000000",
"1101100101111100011010",
"1101100101110110110101",
"1101100101110001001111",
"1101100101101011101001",
"1101100101100110000011",
"1101100101100000011110",
"1101100101011010111000",
"1101100101010101010010",
"1101100101001111101100",
"1101100101001010000111",
"1101100101000100100001",
"1101100100111110111011",
"1101100100111001010101",
"1101100100110011110000",
"1101100100101110001010",
"1101100100101000100100",
"1101100100100010111110",
"1101100100011101011001",
"1101100100010111110011",
"1101100100010010001101",
"1101100100001100100111",
"1101100100000111000010",
"1101100100000001011100",
"1101100011111011110110",
"1101100011110110010000",
"1101100011110000101011",
"1101100011101011000101",
"1101100011100101011111",
"1101100011011111111001",
"1101100011011010010100",
"1101100011010100101110",
"1101100011001111001000",
"1101100011001001100010",
"1101100011000011111101",
"1101100010111110010111",
"1101100010111000110001",
"1101100010110011001011",
"1101100010101101100110",
"1101100010101000000000",
"1101100010100010011010",
"1101100010011100110101",
"1101100010010111001111",
"1101100010010001101001",
"1101100010001100000011",
"1101100010000110011110",
"1101100010000000111000",
"1101100001111011010010",
"1101100001110101101100",
"1101100001110000000111",
"1101100001101010100001",
"1101100001100100111011",
"1101100001011111010101",
"1101100001011001110000",
"1101100001010100001010",
"1101100001001110100100",
"1101100001001000111110",
"1101100001000011011001",
"1101100000111101110011",
"1101100000111000001101",
"1101100000110010100111",
"1101100000101101000010",
"1101100000100111011100",
"1101100000100001110110",
"1101100000011100010000",
"1101100000010110101011",
"1101100000010001000101",
"1101100000001011011111",
"1101100000000101111001",
"1101100000000000010100",
"1101011111111010101110",
"1101011111110101001000",
"1101011111101111100010",
"1101011111101001111101",
"1101011111100100010111",
"1101011111011110110001",
"1101011111011001001011",
"1101011111010011100110",
"1101011111001110000000",
"1101011111001000011010",
"1101011111000010110101",
"1101011110111101001111",
"1101011110110111101001",
"1101011110110010000011",
"1101011110101100011110",
"1101011110100110111000",
"1101011110100001010010",
"1101011110011011101100",
"1101011110010110000111",
"1101011110010000100001",
"1101011110001010111011",
"1101011110000101010101",
"1101011101111111110000",
"1101011101111010001010",
"1101011101110100100100",
"1101011101101110111110",
"1101011101101001011001",
"1101011101100011110011",
"1101011101011110001101",
"1101011101011000100111",
"1101011101010011000010",
"1101011101001101011100",
"1101011101000111110110",
"1101011101000010010000",
"1101011100111100101011",
"1101011100110111000101",
"1101011100110001011111",
"1101011100101011111001",
"1101011100100110010100",
"1101011100100000101110",
"1101011100011011001000",
"1101011100010101100010",
"1101011100001111111101",
"1101011100001010010111",
"1101011100000100110001",
"1101011011111111001011",
"1101011011111001100110",
"1101011011110100000000",
"1101011011101110011010",
"1101011011101000110101",
"1101011011100011001111",
"1101011011011101101001",
"1101011011011000000011",
"1101011011010010011110",
"1101011011001100111000",
"1101011011000111010010",
"1101011011000001101100",
"1101011010111100000111",
"1101011010110110100001",
"1101011010110000111011",
"1101011010101011010101",
"1101011010100101110000",
"1101011010100000001010",
"1101011010011010100100",
"1101011010010100111110",
"1101011010001111011001",
"1101011010001001110011",
"1101011010000100001101",
"1101011001111110100111",
"1101011001111001000010",
"1101011001110011011100",
"1101011001101101110110",
"1101011001101000010000",
"1101011001100010101011",
"1101011001011101000101",
"1101011001010111011111",
"1101011001010001111001",
"1101011001001100010100",
"1101011001000110101110",
"1101011001000001001000",
"1101011000111011100010",
"1101011000110101111101",
"1101011000110000010111",
"1101011000101010110001",
"1101011000100101001011",
"1101011000011111100110",
"1101011000011010000000",
"1101011000010100011010",
"1101011000001110110101",
"1101011000001001001111",
"1101011000000011101001",
"1101010111111110000011",
"1101010111111000011110",
"1101010111110010111000",
"1101010111101101010010",
"1101010111100111101100",
"1101010111100010000111",
"1101010111011100100001",
"1101010111010110111011",
"1101010111010001010101",
"1101010111001011110000",
"1101010111000110001010",
"1101010111000000100100",
"1101010110111010111110",
"1101010110110101011001",
"1101010110101111110011",
"1101010110101010001101",
"1101010110100100100111",
"1101010110011111000010",
"1101010110011001011100",
"1101010110010011110110",
"1101010110001110010000",
"1101010110001000101011",
"1101010110000011000101",
"1101010101111101011111",
"1101010101110111111001",
"1101010101110010010100",
"1101010101101100101110",
"1101010101100111001000",
"1101010101100001100010",
"1101010101011011111101",
"1101010101010110010111",
"1101010101010000110001",
"1101010101001011001011",
"1101010101000101100110",
"1101010101000000000000",
"1101010100111010011010",
"1101010100110100110101",
"1101010100101111001111",
"1101010100101001101001",
"1101010100100100000011",
"1101010100011110011110",
"1101010100011000111000",
"1101010100010011010010",
"1101010100001101101100",
"1101010100001000000111",
"1101010100000010100001",
"1101010011111100111011",
"1101010011110111010101",
"1101010011110001110000",
"1101010011101100001010",
"1101010011100110100100",
"1101010011100000111110",
"1101010011011011011001",
"1101010011010101110011",
"1101010011010000001101",
"1101010011001010100111",
"1101010011000101000010",
"1101010010111111011100",
"1101010010111001110110",
"1101010010110100010000",
"1101010010101110101011",
"1101010010101001000101",
"1101010010100011011111",
"1101010010011101111001",
"1101010010011000010100",
"1101010010010010101110",
"1101010010001101001000",
"1101010010000111100010",
"1101010010000001111101",
"1101010001111100010111",
"1101010001110110110001",
"1101010001110001001011",
"1101010001101011100110",
"1101010001100110000000",
"1101010001100000011010",
"1101010001011010110101",
"1101010001010101001111",
"1101010001001111101001",
"1101010001001010000011",
"1101010001000100011110",
"1101010000111110111000",
"1101010000111001010010",
"1101010000110011101100",
"1101010000101110000111",
"1101010000101000100001",
"1101010000100010111011",
"1101010000011101010101",
"1101010000010111110000",
"1101010000010010001010",
"1101010000001100100100",
"1101010000000110111110",
"1101010000000001011001",
"1101001111111011110011",
"1101001111110110001101",
"1101001111110000100111",
"1101001111101011000010",
"1101001111100101011100",
"1101001111011111110110",
"1101001111011010010000",
"1101001111010100101011",
"1101001111001111000101",
"1101001111001001011111",
"1101001111000011111001",
"1101001110111110010100",
"1101001110111000101110",
"1101001110110011001000",
"1101001110101101100010",
"1101001110100111111101",
"1101001110100010010111",
"1101001110011100110001",
"1101001110010111001011",
"1101001110010001100110",
"1101001110001100000000",
"1101001110000110011010",
"1101001110000000110101",
"1101001101111011001111",
"1101001101110101101001",
"1101001101110000000011",
"1101001101101010011110",
"1101001101100100111000",
"1101001101011111010010",
"1101001101011001101100",
"1101001101010100000111",
"1101001101001110100001",
"1101001101001000111011",
"1101001101000011010101",
"1101001100111101110000",
"1101001100111000001010",
"1101001100110010100100",
"1101001100101100111110",
"1101001100100111011001",
"1101001100100001110011",
"1101001100011100001101",
"1101001100010110100111",
"1101001100010001000010",
"1101001100001011011100",
"1101001100000101110110",
"1101001100000000010000",
"1101001011111010101011",
"1101001011110101000101",
"1101001011101111011111",
"1101001011101001111001",
"1101001011100100010100",
"1101001011011110101110",
"1101001011011001001000",
"1101001011010011100010",
"1101001011001101111101",
"1101001011001000010111",
"1101001011000010110001",
"1101001010111101001011",
"1101001010110111100110",
"1101001010110010000000",
"1101001010101100011010",
"1101001010100110110101",
"1101001010100001001111",
"1101001010011011101001",
"1101001010010110000011",
"1101001010010000011110",
"1101001010001010111000",
"1101001010000101010010",
"1101001001111111101100",
"1101001001111010000111",
"1101001001110100100001",
"1101001001101110111011",
"1101001001101001010101",
"1101001001100011110000",
"1101001001011110001010",
"1101001001011000100100",
"1101001001010010111110",
"1101001001001101011001",
"1101001001000111110011",
"1101001001000010001101",
"1101001000111100100111",
"1101001000110111000010",
"1101001000110001011100",
"1101001000101011110110",
"1101001000100110010000",
"1101001000100000101011",
"1101001000011011000101",
"1101001000010101011111",
"1101001000001111111001",
"1101001000001010010100",
"1101001000000100101110",
"1101000111111111001000",
"1101000111111001100010",
"1101000111110011111101",
"1101000111101110010111",
"1101000111101000110001",
"1101000111100011001011",
"1101000111011101100110",
"1101000111011000000000",
"1101000111010010011010",
"1101000111001100110101",
"1101000111000111001111",
"1101000111000001101001",
"1101000110111100000011",
"1101000110110110011110",
"1101000110110000111000",
"1101000110101011010010",
"1101000110100101101100",
"1101000110100000000111",
"1101000110011010100001",
"1101000110010100111011",
"1101000110001111010101",
"1101000110001001110000",
"1101000110000100001010",
"1101000101111110100100",
"1101000101111000111110",
"1101000101110011011001",
"1101000101101101110011",
"1101000101101000001101",
"1101000101100010100111",
"1101000101011101000010",
"1101000101010111011100",
"1101000101010001110110",
"1101000101001100010000",
"1101000101000110101011",
"1101000101000001000101",
"1101000100111011011111",
"1101000100110101111001",
"1101000100110000010100",
"1101000100101010101110",
"1101000100100101001000",
"1101000100011111100010",
"1101000100011001111101",
"1101000100010100010111",
"1101000100001110110001",
"1101000100001001001011",
"1101000100000011100110",
"1101000011111110000000",
"1101000011111000011010",
"1101000011110010110101",
"1101000011101101001111",
"1101000011100111101001",
"1101000011100010000011",
"1101000011011100011110",
"1101000011010110111000",
"1101000011010001010010",
"1101000011001011101100",
"1101000011000110000111",
"1101000011000000100001",
"1101000010111010111011",
"1101000010110101010101",
"1101000010101111110000",
"1101000010101010001010",
"1101000010100100100100",
"1101000010011110111110",
"1101000010011001011001",
"1101000010010011110011",
"1101000010001110001101",
"1101000010001000100111",
"1101000010000011000010",
"1101000001111101011100",
"1101000001110111110110",
"1101000001110010010000",
"1101000001101100101011",
"1101000001100111000101",
"1101000001100001011111",
"1101000001011011111001",
"1101000001010110010100",
"1101000001010000101110",
"1101000001001011001000",
"1101000001000101100010",
"1101000000111111111101",
"1101000000111010010111",
"1101000000110100110001",
"1101000000101111001011",
"1101000000101001100110",
"1101000000100100000000",
"1101000000011110011010",
"1101000000011000110101",
"1101000000010011001111",
"1101000000001101101001",
"1101000000001000000011",
"1101000000000010011110",
"1100111111111100111000",
"1100111111110111010010",
"1100111111110001101100",
"1100111111101100000111",
"1100111111100110100001",
"1100111111100000111011",
"1100111111011011010101",
"1100111111010101110000",
"1100111111010000001010",
"1100111111001010100100",
"1100111111000100111110",
"1100111110111111011001",
"1100111110111001110011",
"1100111110110100001101",
"1100111110101110100111",
"1100111110101001000010",
"1100111110100011011100",
"1100111110011101110110",
"1100111110011000010000",
"1100111110010010101011",
"1100111110001101000101",
"1100111110000111011111",
"1100111110000001111001",
"1100111101111100010100",
"1100111101110110101110",
"1100111101110001001000",
"1100111101101011100010",
"1100111101100101111101",
"1100111101100000010111",
"1100111101011010110001",
"1100111101010101001011",
"1100111101001111100110",
"1100111101001010000000",
"1100111101000100011010",
"1100111100111110110101",
"1100111100111001001111",
"1100111100110011101001",
"1100111100101110000011",
"1100111100101000011110",
"1100111100100010111000",
"1100111100011101010010",
"1100111100010111101100",
"1100111100010010000111",
"1100111100001100100001",
"1100111100000110111011",
"1100111100000001010101",
"1100111011111011110000",
"1100111011110110001010",
"1100111011110000100100",
"1100111011101010111110",
"1100111011100101011001",
"1100111011011111110011",
"1100111011011010001101",
"1100111011010100100111",
"1100111011001111000010",
"1100111011001001011100",
"1100111011000011110110",
"1100111010111110010000",
"1100111010111000101011",
"1100111010110011000101",
"1100111010101101011111",
"1100111010100111111001",
"1100111010100010010100",
"1100111010011100101110",
"1100111010010111001000",
"1100111010010001100010",
"1100111010001011111101",
"1100111010000110010111",
"1100111010000000110001",
"1100111001111011001011",
"1100111001110101100110",
"1100111001110000000000",
"1100111001101010011010",
"1100111001100100110101",
"1100111001011111001111",
"1100111001011001101001",
"1100111001010100000011",
"1100111001001110011110",
"1100111001001000111000",
"1100111001000011010010",
"1100111000111101101100",
"1100111000111000000111",
"1100111000110010100001",
"1100111000101100111011",
"1100111000100111010101",
"1100111000100001110000",
"1100111000011100001010",
"1100111000010110100100",
"1100111000010000111110",
"1100111000001011011001",
"1100111000000101110011",
"1100111000000000001101",
"1100110111111010100111",
"1100110111110101000010",
"1100110111101111011100",
"1100110111101001110110",
"1100110111100100010000",
"1100110111011110101011",
"1100110111011001000101",
"1100110111010011011111",
"1100110111001101111001",
"1100110111001000010100",
"1100110111000010101110",
"1100110110111101001000",
"1100110110110111100010",
"1100110110110001111101",
"1100110110101100010111",
"1100110110100110110001",
"1100110110100001001011",
"1100110110011011100110",
"1100110110010110000000",
"1100110110010000011010",
"1100110110001010110101",
"1100110110000101001111",
"1100110101111111101001",
"1100110101111010000011",
"1100110101110100011110",
"1100110101101110111000",
"1100110101101001010010",
"1100110101100011101100",
"1100110101011110000111",
"1100110101011000100001",
"1100110101010010111011",
"1100110101001101010101",
"1100110101000111110000",
"1100110101000010001010",
"1100110100111100100100",
"1100110100110110111110",
"1100110100110001011001",
"1100110100101011110011",
"1100110100100110001101",
"1100110100100000100111",
"1100110100011011000010",
"1100110100010101011100",
"1100110100001111110110",
"1100110100001010010000",
"1100110100000100101011",
"1100110011111111000101",
"1100110011111001011111",
"1100110011110011111001",
"1100110011101110010100",
"1100110011101000101110",
"1100110011100011001000",
"1100110011011101100010",
"1100110011010111111101",
"1100110011010010010111",
"1100110011001100110001",
"1100110011000111001011",
"1100110011000001100110",
"1100110010111100000000",
"1100110010110110011010",
"1100110010110000110101",
"1100110010101011001111",
"1100110010100101101001",
"1100110010100000000011",
"1100110010011010011110",
"1100110010010100111000",
"1100110010001111010010",
"1100110010001001101100",
"1100110010000100000111",
"1100110001111110100001",
"1100110001111000111011",
"1100110001110011010101",
"1100110001101101110000",
"1100110001101000001010",
"1100110001100010100100",
"1100110001011100111110",
"1100110001010111011001",
"1100110001010001110011",
"1100110001001100001101",
"1100110001000110100111",
"1100110001000001000010",
"1100110000111011011100",
"1100110000110101110110",
"1100110000110000010000",
"1100110000101010101011",
"1100110000100101000101",
"1100110000011111011111",
"1100110000011001111001",
"1100110000010100010100",
"1100110000001110101110",
"1100110000001001001000",
"1100110000000011100010",
"1100101111111101111101",
"1100101111111000010111",
"1100101111110010110001",
"1100101111101101001011",
"1100101111100111100110",
"1100101111100010000000",
"1100101111011100011010",
"1100101111010110110101",
"1100101111010001001111",
"1100101111001011101001",
"1100101111000110000011",
"1100101111000000011110",
"1100101110111010111000",
"1100101110110101010010",
"1100101110101111101100",
"1100101110101010000111",
"1100101110100100100001",
"1100101110011110111011",
"1100101110011001010101",
"1100101110010011110000",
"1100101110001110001010",
"1100101110001000100100",
"1100101110000010111110",
"1100101101111101011001",
"1100101101110111110011",
"1100101101110010001101",
"1100101101101100100111",
"1100101101100111000010",
"1100101101100001011100",
"1100101101011011110110",
"1100101101010110010000",
"1100101101010000101011",
"1100101101001011000101",
"1100101101000101011111",
"1100101100111111111001",
"1100101100111010010100",
"1100101100110100101110",
"1100101100101111001000",
"1100101100101001100010",
"1100101100100011111101",
"1100101100011110010111",
"1100101100011000110001",
"1100101100010011001011",
"1100101100001101100110",
"1100101100001000000000",
"1100101100000010011010",
"1100101011111100110101",
"1100101011110111001111",
"1100101011110001101001",
"1100101011101100000011",
"1100101011100110011110",
"1100101011100000111000",
"1100101011011011010010",
"1100101011010101101100",
"1100101011010000000111",
"1100101011001010100001",
"1100101011000100111011",
"1100101010111111010101",
"1100101010111001110000",
"1100101010110100001010",
"1100101010101110100100",
"1100101010101000111110",
"1100101010100011011001",
"1100101010011101110011",
"1100101010011000001101",
"1100101010010010100111",
"1100101010001101000010",
"1100101010000111011100",
"1100101010000001110110",
"1100101001111100010000",
"1100101001110110101011",
"1100101001110001000101",
"1100101001101011011111",
"1100101001100101111001",
"1100101001100000010100",
"1100101001011010101110",
"1100101001010101001000",
"1100101001001111100010",
"1100101001001001111101",
"1100101001000100010111",
"1100101000111110110001",
"1100101000111001001011",
"1100101000110011100110",
"1100101000101110000000",
"1100101000101000011010",
"1100101000100010110101",
"1100101000011101001111",
"1100101000010111101001",
"1100101000010010000011",
"1100101000001100011110",
"1100101000000110111000",
"1100101000000001010010",
"1100100111111011101100",
"1100100111110110000111",
"1100100111110000100001",
"1100100111101010111011",
"1100100111100101010101",
"1100100111011111110000",
"1100100111011010001010",
"1100100111010100100100",
"1100100111001110111110",
"1100100111001001011001",
"1100100111000011110011",
"1100100110111110001101",
"1100100110111000100111",
"1100100110110011000010",
"1100100110101101011100",
"1100100110100111110110",
"1100100110100010010000",
"1100100110011100101011",
"1100100110010111000101",
"1100100110010001011111",
"1100100110001011111001",
"1100100110000110010100",
"1100100110000000101110",
"1100100101111011001000",
"1100100101110101100010",
"1100100101101111111101",
"1100100101101010010111",
"1100100101100100110001",
"1100100101011111001011",
"1100100101011001100110",
"1100100101010100000000",
"1100100101001110011010",
"1100100101001000110101",
"1100100101000011001111",
"1100100100111101101001",
"1100100100111000000011",
"1100100100110010011110",
"1100100100101100111000",
"1100100100100111010010",
"1100100100100001101100",
"1100100100011100000111",
"1100100100010110100001",
"1100100100010000111011",
"1100100100001011010101",
"1100100100000101110000",
"1100100100000000001010",
"1100100011111010100100",
"1100100011110100111110",
"1100100011101111011001",
"1100100011101001110011",
"1100100011100100001101",
"1100100011011110100111",
"1100100011011001000010",
"1100100011010011011100",
"1100100011001101110110",
"1100100011001000010000",
"1100100011000010101011",
"1100100010111101000101",
"1100100010110111011111",
"1100100010110001111001",
"1100100010101100010100",
"1100100010100110101110",
"1100100010100001001000",
"1100100010011011100010",
"1100100010010101111101",
"1100100010010000010111",
"1100100010001010110001",
"1100100010000101001011",
"1100100001111111100110",
"1100100001111010000000",
"1100100001110100011010",
"1100100001101110110101",
"1100100001101001001111",
"1100100001100011101001",
"1100100001011110000011",
"1100100001011000011110",
"1100100001010010111000",
"1100100001001101010010",
"1100100001000111101100",
"1100100001000010000111",
"1100100000111100100001",
"1100100000110110111011",
"1100100000110001010101",
"1100100000101011110000",
"1100100000100110001010",
"1100100000100000100100",
"1100100000011010111110",
"1100100000010101011001",
"1100100000001111110011",
"1100100000001010001101",
"1100100000000100100111",
"1100011111111111000010",
"1100011111111001011100",
"1100011111110011110110",
"1100011111101110010000",
"1100011111101000101011",
"1100011111100011000101",
"1100011111011101011111",
"1100011111010111111001",
"1100011111010010010100",
"1100011111001100101110",
"1100011111000111001000",
"1100011111000001100010",
"1100011110111011111101",
"1100011110110110010111",
"1100011110110000110001",
"1100011110101011001011",
"1100011110100101100110",
"1100011110100000000000",
"1100011110011010011010",
"1100011110010100110101",
"1100011110001111001111",
"1100011110001001101001",
"1100011110000100000011",
"1100011101111110011110",
"1100011101111000111000",
"1100011101110011010010",
"1100011101101101101100",
"1100011101101000000111",
"1100011101100010100001",
"1100011101011100111011",
"1100011101010111010101",
"1100011101010001110000",
"1100011101001100001010",
"1100011101000110100100",
"1100011101000000111110",
"1100011100111011011001",
"1100011100110101110011",
"1100011100110000001101",
"1100011100101010100111",
"1100011100100101000010",
"1100011100011111011100",
"1100011100011001110110",
"1100011100010100010000",
"1100011100001110101011",
"1100011100001001000101",
"1100011100000011011111",
"1100011011111101111001",
"1100011011111000010100",
"1100011011110010101110",
"1100011011101101001000",
"1100011011100111100010",
"1100011011100001111101",
"1100011011011100010111",
"1100011011010110110001",
"1100011011010001001011",
"1100011011001011100110",
"1100011011000110000000",
"1100011011000000011010",
"1100011010111010110101",
"1100011010110101001111",
"1100011010101111101001",
"1100011010101010000011",
"1100011010100100011110",
"1100011010011110111000",
"1100011010011001010010",
"1100011010010011101100",
"1100011010001110000111",
"1100011010001000100001",
"1100011010000010111011",
"1100011001111101010101",
"1100011001110111110000",
"1100011001110010001010",
"1100011001101100100100",
"1100011001100110111110",
"1100011001100001011001",
"1100011001011011110011",
"1100011001010110001101",
"1100011001010000100111",
"1100011001001011000010",
"1100011001000101011100",
"1100011000111111110110",
"1100011000111010010000",
"1100011000110100101011",
"1100011000101111000101",
"1100011000101001011111",
"1100011000100011111001",
"1100011000011110010100",
"1100011000011000101110",
"1100011000010011001000",
"1100011000001101100010",
"1100011000000111111101",
"1100011000000010010111",
"1100010111111100110001",
"1100010111110111001011",
"1100010111110001100110",
"1100010111101100000000",
"1100010111100110011010",
"1100010111100000110101",
"1100010111011011001111",
"1100010111010101101001",
"1100010111010000000011",
"1100010111001010011110",
"1100010111000100111000",
"1100010110111111010010",
"1100010110111001101100",
"1100010110110100000111",
"1100010110101110100001",
"1100010110101000111011",
"1100010110100011010101",
"1100010110011101110000",
"1100010110011000001010",
"1100010110010010100100",
"1100010110001100111110",
"1100010110000111011001",
"1100010110000001110011",
"1100010101111100001101",
"1100010101110110100111",
"1100010101110001000010",
"1100010101101011011100",
"1100010101100101110110",
"1100010101100000010000",
"1100010101011010101011",
"1100010101010101000101",
"1100010101001111011111",
"1100010101001001111001",
"1100010101000100010100",
"1100010100111110101110",
"1100010100111001001000",
"1100010100110011100010"
    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
				
				mem_out_reg(21 downto 0) <= mem_out_next(21 downto 0);
  
     --       if we = '1' then
     --           mem(to_integer(unsigned(addr))) <= d_in;  -- Write operation
     --      end if;
        end if;
    end process;
	 
		mem_out_next <= mem(to_integer(unsigned(addr)));      -- Read operation
		d_out(21 downto 0) <= mem_out_reg(21 downto 0); 
	 
	 
	 
end rtl;