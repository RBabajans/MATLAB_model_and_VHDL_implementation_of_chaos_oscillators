library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Exponent_memory is
    Port (
        clk      : in  STD_LOGIC;  -- Clock signal
        we       : in  STD_LOGIC;  -- Write Enable
        addr     : in  STD_LOGIC_VECTOR(11 downto 0); -- 12-bit Address space
        d_in      : in  STD_LOGIC_VECTOR(21 downto 0); -- Data input (22-bit)
        d_out     : out STD_LOGIC_VECTOR(21 downto 0)  -- Data output (22-bit)
    );
end Exponent_memory;

architecture rtl of Exponent_memory is

	 signal mem_out_reg, mem_out_next : STD_LOGIC_VECTOR(21 downto 0) := (others => '0');


    type Heaviside_Array is array (0 to 4095) of STD_LOGIC_VECTOR(21 downto 0);  -- Memory array
    signal mem : Heaviside_Array := (
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011101",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011100",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011011",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011010",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011001",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001011000",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010111",
		"0010000011100001010110",
		"0010000011100001010110",
		"0010000011100001010110",
		"0010000011100001010110",
		"0010000011100001010110",
		"0010000011100001010110",
		"0010000011100001010110",
		"0010000011100001010110",
		"0010000011100001010110",
		"0010000011100001010101",
		"0010000011100001010101",
		"0010000011100001010101",
		"0010000011100001010101",
		"0010000011100001010101",
		"0010000011100001010101",
		"0010000011100001010101",
		"0010000011100001010101",
		"0010000011100001010101",
		"0010000011100001010100",
		"0010000011100001010100",
		"0010000011100001010100",
		"0010000011100001010100",
		"0010000011100001010100",
		"0010000011100001010100",
		"0010000011100001010100",
		"0010000011100001010011",
		"0010000011100001010011",
		"0010000011100001010011",
		"0010000011100001010011",
		"0010000011100001010011",
		"0010000011100001010011",
		"0010000011100001010010",
		"0010000011100001010010",
		"0010000011100001010010",
		"0010000011100001010010",
		"0010000011100001010010",
		"0010000011100001010010",
		"0010000011100001010001",
		"0010000011100001010001",
		"0010000011100001010001",
		"0010000011100001010001",
		"0010000011100001010001",
		"0010000011100001010001",
		"0010000011100001010000",
		"0010000011100001010000",
		"0010000011100001010000",
		"0010000011100001010000",
		"0010000011100001010000",
		"0010000011100001001111",
		"0010000011100001001111",
		"0010000011100001001111",
		"0010000011100001001111",
		"0010000011100001001111",
		"0010000011100001001110",
		"0010000011100001001110",
		"0010000011100001001110",
		"0010000011100001001110",
		"0010000011100001001101",
		"0010000011100001001101",
		"0010000011100001001101",
		"0010000011100001001101",
		"0010000011100001001100",
		"0010000011100001001100",
		"0010000011100001001100",
		"0010000011100001001100",
		"0010000011100001001011",
		"0010000011100001001011",
		"0010000011100001001011",
		"0010000011100001001010",
		"0010000011100001001010",
		"0010000011100001001010",
		"0010000011100001001010",
		"0010000011100001001001",
		"0010000011100001001001",
		"0010000011100001001001",
		"0010000011100001001000",
		"0010000011100001001000",
		"0010000011100001001000",
		"0010000011100001000111",
		"0010000011100001000111",
		"0010000011100001000111",
		"0010000011100001000110",
		"0010000011100001000110",
		"0010000011100001000110",
		"0010000011100001000101",
		"0010000011100001000101",
		"0010000011100001000101",
		"0010000011100001000100",
		"0010000011100001000100",
		"0010000011100001000011",
		"0010000011100001000011",
		"0010000011100001000011",
		"0010000011100001000010",
		"0010000011100001000010",
		"0010000011100001000001",
		"0010000011100001000001",
		"0010000011100001000000",
		"0010000011100001000000",
		"0010000011100001000000",
		"0010000011100000111111",
		"0010000011100000111111",
		"0010000011100000111110",
		"0010000011100000111110",
		"0010000011100000111101",
		"0010000011100000111101",
		"0010000011100000111100",
		"0010000011100000111100",
		"0010000011100000111011",
		"0010000011100000111011",
		"0010000011100000111010",
		"0010000011100000111010",
		"0010000011100000111001",
		"0010000011100000111000",
		"0010000011100000111000",
		"0010000011100000110111",
		"0010000011100000110111",
		"0010000011100000110110",
		"0010000011100000110101",
		"0010000011100000110101",
		"0010000011100000110100",
		"0010000011100000110100",
		"0010000011100000110011",
		"0010000011100000110010",
		"0010000011100000110010",
		"0010000011100000110001",
		"0010000011100000110000",
		"0010000011100000101111",
		"0010000011100000101111",
		"0010000011100000101110",
		"0010000011100000101101",
		"0010000011100000101101",
		"0010000011100000101100",
		"0010000011100000101011",
		"0010000011100000101010",
		"0010000011100000101001",
		"0010000011100000101001",
		"0010000011100000101000",
		"0010000011100000100111",
		"0010000011100000100110",
		"0010000011100000100101",
		"0010000011100000100100",
		"0010000011100000100100",
		"0010000011100000100011",
		"0010000011100000100010",
		"0010000011100000100001",
		"0010000011100000100000",
		"0010000011100000011111",
		"0010000011100000011110",
		"0010000011100000011101",
		"0010000011100000011100",
		"0010000011100000011011",
		"0010000011100000011010",
		"0010000011100000011001",
		"0010000011100000011000",
		"0010000011100000010111",
		"0010000011100000010110",
		"0010000011100000010100",
		"0010000011100000010011",
		"0010000011100000010010",
		"0010000011100000010001",
		"0010000011100000010000",
		"0010000011100000001111",
		"0010000011100000001101",
		"0010000011100000001100",
		"0010000011100000001011",
		"0010000011100000001010",
		"0010000011100000001000",
		"0010000011100000000111",
		"0010000011100000000110",
		"0010000011100000000100",
		"0010000011100000000011",
		"0010000011100000000001",
		"0010000011100000000000",
		"0010000011011111111110",
		"0010000011011111111101",
		"0010000011011111111011",
		"0010000011011111111010",
		"0010000011011111111000",
		"0010000011011111110111",
		"0010000011011111110101",
		"0010000011011111110100",
		"0010000011011111110010",
		"0010000011011111110000",
		"0010000011011111101110",
		"0010000011011111101101",
		"0010000011011111101011",
		"0010000011011111101001",
		"0010000011011111100111",
		"0010000011011111100110",
		"0010000011011111100100",
		"0010000011011111100010",
		"0010000011011111100000",
		"0010000011011111011110",
		"0010000011011111011100",
		"0010000011011111011010",
		"0010000011011111011000",
		"0010000011011111010110",
		"0010000011011111010100",
		"0010000011011111010001",
		"0010000011011111001111",
		"0010000011011111001101",
		"0010000011011111001011",
		"0010000011011111001000",
		"0010000011011111000110",
		"0010000011011111000100",
		"0010000011011111000001",
		"0010000011011110111111",
		"0010000011011110111100",
		"0010000011011110111010",
		"0010000011011110110111",
		"0010000011011110110101",
		"0010000011011110110010",
		"0010000011011110101111",
		"0010000011011110101101",
		"0010000011011110101010",
		"0010000011011110100111",
		"0010000011011110100100",
		"0010000011011110100001",
		"0010000011011110011110",
		"0010000011011110011011",
		"0010000011011110011000",
		"0010000011011110010101",
		"0010000011011110010010",
		"0010000011011110001111",
		"0010000011011110001100",
		"0010000011011110001000",
		"0010000011011110000101",
		"0010000011011110000001",
		"0010000011011101111110",
		"0010000011011101111011",
		"0010000011011101110111",
		"0010000011011101110011",
		"0010000011011101110000",
		"0010000011011101101100",
		"0010000011011101101000",
		"0010000011011101100100",
		"0010000011011101100000",
		"0010000011011101011100",
		"0010000011011101011000",
		"0010000011011101010100",
		"0010000011011101010000",
		"0010000011011101001100",
		"0010000011011101001000",
		"0010000011011101000011",
		"0010000011011100111111",
		"0010000011011100111010",
		"0010000011011100110110",
		"0010000011011100110001",
		"0010000011011100101100",
		"0010000011011100101000",
		"0010000011011100100011",
		"0010000011011100011110",
		"0010000011011100011001",
		"0010000011011100010100",
		"0010000011011100001110",
		"0010000011011100001001",
		"0010000011011100000100",
		"0010000011011011111110",
		"0010000011011011111001",
		"0010000011011011110011",
		"0010000011011011101110",
		"0010000011011011101000",
		"0010000011011011100010",
		"0010000011011011011100",
		"0010000011011011010110",
		"0010000011011011010000",
		"0010000011011011001001",
		"0010000011011011000011",
		"0010000011011010111101",
		"0010000011011010110110",
		"0010000011011010101111",
		"0010000011011010101001",
		"0010000011011010100010",
		"0010000011011010011011",
		"0010000011011010010100",
		"0010000011011010001101",
		"0010000011011010000101",
		"0010000011011001111110",
		"0010000011011001110110",
		"0010000011011001101111",
		"0010000011011001100111",
		"0010000011011001011111",
		"0010000011011001010111",
		"0010000011011001001111",
		"0010000011011001000110",
		"0010000011011000111110",
		"0010000011011000110110",
		"0010000011011000101101",
		"0010000011011000100100",
		"0010000011011000011011",
		"0010000011011000010010",
		"0010000011011000001001",
		"0010000011010111111111",
		"0010000011010111110110",
		"0010000011010111101100",
		"0010000011010111100010",
		"0010000011010111011000",
		"0010000011010111001110",
		"0010000011010111000100",
		"0010000011010110111001",
		"0010000011010110101111",
		"0010000011010110100100",
		"0010000011010110011001",
		"0010000011010110001110",
		"0010000011010110000010",
		"0010000011010101110111",
		"0010000011010101101011",
		"0010000011010101011111",
		"0010000011010101010011",
		"0010000011010101000111",
		"0010000011010100111011",
		"0010000011010100101110",
		"0010000011010100100001",
		"0010000011010100010100",
		"0010000011010100000111",
		"0010000011010011111010",
		"0010000011010011101100",
		"0010000011010011011110",
		"0010000011010011010000",
		"0010000011010011000010",
		"0010000011010010110011",
		"0010000011010010100100",
		"0010000011010010010101",
		"0010000011010010000110",
		"0010000011010001110111",
		"0010000011010001100111",
		"0010000011010001010111",
		"0010000011010001000111",
		"0010000011010000110110",
		"0010000011010000100101",
		"0010000011010000010100",
		"0010000011010000000011",
		"0010000011001111110010",
		"0010000011001111100000",
		"0010000011001111001110",
		"0010000011001110111011",
		"0010000011001110101001",
		"0010000011001110010110",
		"0010000011001110000011",
		"0010000011001101101111",
		"0010000011001101011011",
		"0010000011001101000111",
		"0010000011001100110010",
		"0010000011001100011110",
		"0010000011001100001000",
		"0010000011001011110011",
		"0010000011001011011101",
		"0010000011001011000111",
		"0010000011001010110000",
		"0010000011001010011010",
		"0010000011001010000010",
		"0010000011001001101011",
		"0010000011001001010011",
		"0010000011001000111010",
		"0010000011001000100010",
		"0010000011001000001001",
		"0010000011000111101111",
		"0010000011000111010101",
		"0010000011000110111011",
		"0010000011000110100000",
		"0010000011000110000101",
		"0010000011000101101001",
		"0010000011000101001101",
		"0010000011000100110001",
		"0010000011000100010100",
		"0010000011000011110111",
		"0010000011000011011001",
		"0010000011000010111010",
		"0010000011000010011100",
		"0010000011000001111100",
		"0010000011000001011101",
		"0010000011000000111100",
		"0010000011000000011100",
		"0010000010111111111010",
		"0010000010111111011001",
		"0010000010111110110110",
		"0010000010111110010011",
		"0010000010111101110000",
		"0010000010111101001100",
		"0010000010111100100111",
		"0010000010111100000010",
		"0010000010111011011101",
		"0010000010111010110110",
		"0010000010111010001111",
		"0010000010111001101000",
		"0010000010111001000000",
		"0010000010111000010111",
		"0010000010110111101110",
		"0010000010110111000011",
		"0010000010110110011001",
		"0010000010110101101101",
		"0010000010110101000001",
		"0010000010110100010100",
		"0010000010110011100111",
		"0010000010110010111001",
		"0010000010110010001010",
		"0010000010110001011010",
		"0010000010110000101010",
		"0010000010101111111001",
		"0010000010101111000111",
		"0010000010101110010100",
		"0010000010101101100000",
		"0010000010101100101100",
		"0010000010101011110111",
		"0010000010101011000001",
		"0010000010101010001010",
		"0010000010101001010010",
		"0010000010101000011010",
		"0010000010100111100000",
		"0010000010100110100110",
		"0010000010100101101010",
		"0010000010100100101110",
		"0010000010100011110001",
		"0010000010100010110011",
		"0010000010100001110100",
		"0010000010100000110011",
		"0010000010011111110010",
		"0010000010011110110000",
		"0010000010011101101101",
		"0010000010011100101001",
		"0010000010011011100011",
		"0010000010011010011101",
		"0010000010011001010101",
		"0010000010011000001101",
		"0010000010010111000011",
		"0010000010010101111000",
		"0010000010010100101100",
		"0010000010010011011110",
		"0010000010010010010000",
		"0010000010010001000000",
		"0010000010001111101111",
		"0010000010001110011100",
		"0010000010001101001001",
		"0010000010001011110100",
		"0010000010001010011101",
		"0010000010001001000110",
		"0010000010000111101101",
		"0010000010000110010010",
		"0010000010000100110110",
		"0010000010000011011001",
		"0010000010000001111010",
		"0010000010000000011010",
		"0010000001111110111000",
		"0010000001111101010101",
		"0010000001111011110000",
		"0010000001111010001001",
		"0010000001111000100001",
		"0010000001110110111000",
		"0010000001110101001100",
		"0010000001110011011111",
		"0010000001110001110000",
		"0010000001110000000000",
		"0010000001101110001101",
		"0010000001101100011001",
		"0010000001101010100011",
		"0010000001101000101011",
		"0010000001100110110010",
		"0010000001100100110110",
		"0010000001100010111000",
		"0010000001100000111001",
		"0010000001011110110111",
		"0010000001011100110100",
		"0010000001011010101110",
		"0010000001011000100110",
		"0010000001010110011100",
		"0010000001010100010000",
		"0010000001010010000010",
		"0010000001001111110001",
		"0010000001001101011110",
		"0010000001001011001001",
		"0010000001001000110010",
		"0010000001000110011000",
		"0010000001000011111100",
		"0010000001000001011101",
		"0010000000111110111100",
		"0010000000111100011000",
		"0010000000111001110001",
		"0010000000110111001000",
		"0010000000110100011101",
		"0010000000110001101110",
		"0010000000101110111101",
		"0010000000101100001001",
		"0010000000101001010011",
		"0010000000100110011001",
		"0010000000100011011101",
		"0010000000100000011101",
		"0010000000011101011011",
		"0010000000011010010101",
		"0010000000010111001100",
		"0010000000010100000000",
		"0010000000010000110001",
		"0010000000001101011111",
		"0010000000001010001001",
		"0010000000000110110000",
		"0010000000000011010100",
		"0001111111111111110100",
		"0001111111111100010001",
		"0001111111111000101010",
		"0001111111110100111111",
		"0001111111110001010001",
		"0001111111101101011111",
		"0001111111101001101001",
		"0001111111100101101111",
		"0001111111100001110001",
		"0001111111011101110000",
		"0001111111011001101010",
		"0001111111010101100000",
		"0001111111010001010010",
		"0001111111001101000000",
		"0001111111001000101001",
		"0001111111000100001110",
		"0001111110111111101111",
		"0001111110111011001011",
		"0001111110110110100010",
		"0001111110110001110101",
		"0001111110101101000011",
		"0001111110101000001100",
		"0001111110100011010000",
		"0001111110011110010000",
		"0001111110011001001010",
		"0001111110010011111111",
		"0001111110001110101111",
		"0001111110001001011010",
		"0001111110000011111111",
		"0001111101111110011111",
		"0001111101111000111001",
		"0001111101110011001101",
		"0001111101101101011100",
		"0001111101100111100101",
		"0001111101100001101001",
		"0001111101011011100110",
		"0001111101010101011101",
		"0001111101001111001110",
		"0001111101001000111000",
		"0001111101000010011100",
		"0001111100111011111010",
		"0001111100110101010001",
		"0001111100101110100010",
		"0001111100100111101011",
		"0001111100100000101110",
		"0001111100011001101010",
		"0001111100010010011111",
		"0001111100001011001100",
		"0001111100000011110010",
		"0001111011111100010001",
		"0001111011110100101000",
		"0001111011101100110111",
		"0001111011100100111110",
		"0001111011011100111110",
		"0001111011010100110101",
		"0001111011001100100101",
		"0001111011000100001100",
		"0001111010111011101010",
		"0001111010110011000000",
		"0001111010101010001101",
		"0001111010100001010001",
		"0001111010011000001101",
		"0001111010001110111111",
		"0001111010000101101000",
		"0001111001111100000111",
		"0001111001110010011101",
		"0001111001101000101001",
		"0001111001011110101011",
		"0001111001010100100100",
		"0001111001001010010010",
		"0001111000111111110101",
		"0001111000110101001110",
		"0001111000101010011101",
		"0001111000011111100000",
		"0001111000010100011001",
		"0001111000001001000110",
		"0001110111111101101000",
		"0001110111110001111110",
		"0001110111100110001001",
		"0001110111011010001000",
		"0001110111001101111010",
		"0001110111000001100000",
		"0001110110110100111010",
		"0001110110101000000111",
		"0001110110011011001000",
		"0001110110001101111011",
		"0001110110000000100000",
		"0001110101110010111001",
		"0001110101100101000011",
		"0001110101010111000000",
		"0001110101001000101110",
		"0001110100111010001110",
		"0001110100101011100000",
		"0001110100011100100010",
		"0001110100001101010110",
		"0001110011111101111010",
		"0001110011101110001111",
		"0001110011011110010011",
		"0001110011001110001000",
		"0001110010111101101101",
		"0001110010101101000001",
		"0001110010011100000100",
		"0001110010001010110110",
		"0001110001111001010110",
		"0001110001100111100101",
		"0001110001010101100011",
		"0001110001000011001110",
		"0001110000110000100110",
		"0001110000011101101100",
		"0001110000001010011110",
		"0001101111110110111110",
		"0001101111100011001001",
		"0001101111001111000001",
		"0001101110111010100100",
		"0001101110100101110011",
		"0001101110010000101101",
		"0001101101111011010010",
		"0001101101100101100001",
		"0001101101001111011010",
		"0001101100111000111100",
		"0001101100100010001000",
		"0001101100001010111110",
		"0001101011110011011011",
		"0001101011011011100001",
		"0001101011000011001111",
		"0001101010101010100101",
		"0001101010010001100001",
		"0001101001111000000101",
		"0001101001011110001111",
		"0001101001000011111110",
		"0001101000101001010011",
		"0001101000001110001110",
		"0001100111110010101101",
		"0001100111010110110000",
		"0001100110111010010111",
		"0001100110011101100010",
		"0001100110000000001111",
		"0001100101100010011111",
		"0001100101000100010001",
		"0001100100100101100101",
		"0001100100000110011001",
		"0001100011100110101111",
		"0001100011000110100100",
		"0001100010100101111001",
		"0001100010000100101100",
		"0001100001100010111111",
		"0001100001000000101111",
		"0001100000011101111101",
		"0001011111111010101000",
		"0001011111010110101111",
		"0001011110110010010011",
		"0001011110001101010001",
		"0001011101100111101010",
		"0001011101000001011101",
		"0001011100011010101010",
		"0001011011110011001111",
		"0001011011001011001101",
		"0001011010100010100011",
		"0001011001111001001111",
		"0001011001001111010010",
		"0001011000100100101011",
		"0001010111111001011000",
		"0001010111001101011010",
		"0001010110100000110000",
		"0001010101110011011001",
		"0001010101000101010100",
		"0001010100010110100000",
		"0001010011100110111101",
		"0001010010110110101011",
		"0001010010000101101000",
		"0001010001010011110011",
		"0001010000100001001100",
		"0001001111101101110010",
		"0001001110111001100100",
		"0001001110000100100010",
		"0001001101001110101010",
		"0001001100010111111100",
		"0001001011100000010111",
		"0001001010100111111010",
		"0001001001101110100100",
		"0001001000110100010100",
		"0001000111111001001001",
		"0001000110111101000011",
		"0001000110000000000000",
		"0001000101000010000000",
		"0001000100000011000001",
		"0001000011000011000010",
		"0001000010000010000100",
		"0001000001000000000011",
		"0000111111111101000000",
		"0000111110111000111010",
		"0000111101110011101111",
		"0000111100101101011110",
		"0000111011100110000111",
		"0000111010011101100111",
		"0000111001010011111111",
		"0000111000001001001100",
		"0000110110111101001110",
		"0000110101110000000011",
		"0000110100100001101010",
		"0000110011010010000011",
		"0000110010000001001011",
		"0000110000101111000010",
		"0000101111011011100110",
		"0000101110000110110110",
		"0000101100110000110000",
		"0000101011011001010100",
		"0000101010000000100000",
		"0000101000100110010010",
		"0000100111001010101001",
		"0000100101101101100011",
		"0000100100001111000000",
		"0000100010101110111110",
		"0000100001001101011011",
		"0000011111101010010110",
		"0000011110000101101100",
		"0000011100011111011101",
		"0000011010110111101000",
		"0000011001001110001001",
		"0000010111100011000001",
		"0000010101110110001100",
		"0000010100000111101001",
		"0000010010010111011000",
		"0000010000100101010101",
		"0000001110110001011111",
		"0000001100111011110100",
		"0000001011000100010011",
		"0000001001001010111001",
		"0000000111001111100101",
		"0000000101010010010101",
		"0000000011010011000110",
		"0000000001010001110111",
		"1111111111001110100110",
		"1111111101001001010001",
		"1111111011000001110101",
		"1111111000111000010001",
		"1111110110101100100010",
		"1111110100011110100111",
		"1111110010001110011100",
		"1111101111111100000000",
		"1111101101100111010000",
		"1111101011010000001011",
		"1111101000110110101101",
		"1111100110011010110100",
		"1111100011111100011111",
		"1111100001011011101010",
		"1111011110111000010010",
		"1111011100010010010110",
		"1111011001101001110011",
		"1111010110111110100110",
		"1111010100010000101101",
		"1111010001100000000100",
		"1111001110101100101001",
		"1111001011110110011001",
		"1111001000111101010010",
		"1111000110000001010000",
		"1111000011000010010000",
		"1111000000000000010001",
		"1110111100111011001101",
		"1110111001110011000011",
		"1110110110100111101111",
		"1110110011011001001111",
		"1110110000000111011110",
		"1110101100110010011001",
		"1110101001011001111110",
		"1110100101111110001001",
		"1110100010011110110111",
		"1110011110111100000011",
		"1110011011010101101011",
		"1110010111101011101010",
		"1110010011111101111110",
		"1110010000001100100010",
		"1110001100010111010011",
		"1110001000011110001100",
		"1110000100100001001011",
		"1110000000100000001011",
		"1101111100011011000111",
		"1101111000010001111100",
		"1101110100000100100111",
		"1101101111110011000001",
		"1101101011011101001000",
		"1101100111000010110111",
		"1101100010100100001010",
		"1101011110000000111011",
		"1101011001011001000111",
		"1101010100101100101001",
		"1101001111111011011100",
		"1101001011000101011011",
		"1101000110001010100010",
		"1101000001001010101100",
		"1100111100000101110011",
		"1100110110111011110011",
		"1100110001101100100110",
		"1100101100011000000111",
		"1100100110111110010010",
		"1100100001011110111111",
		"1100011011111010001011",
		"1100010110001111101111",
		"1100010000011111100101",
		"1100001010101001101001",
		"1100000100101101110100",
		"1011111110101100000000",
		"1011111000100100000111",
		"1011110010010110000011",
		"1011101100000001101110",
		"1011100101100111000010",
		"1011011111000101110111",
		"1011011000011110001000",
		"1011010001101111101110",
		"1011001010111010100010",
		"1011000011111110011110",
		"1010111100111011011010",
		"1010110101110001010000",
		"1010101110011111110111",
		"1010100111000111001010",
		"1010011111100111000000",
		"1010010111111111010011",
		"1010010000001111111001",
		"1010001000011000101101",
		"1010000000011001100101",
		"1001111000010010011010",
		"1001110000000011000100",
		"1001100111101011011011",
		"1001011111001011010110",
		"1001010110100010101100",
		"1001001101110001010101",
		"1001000100110111001001",
		"1000111011110011111110",
		"1000110010100111101011",
		"1000101001010010000111",
		"1000011111110011001001",
		"1000010110001010100111",
		"1000001100011000011000",
		"1000000010011100010010",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000",
		"1000000000000000000000"
    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
				
				mem_out_reg(21 downto 0) <= mem_out_next(21 downto 0);
  
        end if;
    end process;
	 
		mem_out_next <= mem(to_integer(unsigned(addr)));      -- Read operation
		d_out(21 downto 0) <= mem_out_reg(21 downto 0); 
	 
	 
	 
end rtl;